  LIBRARY ieee; USE ieee.std_logic_1164.ALL; LIBRARY XilinxCoreLib; ENTITY Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692 IS   PORT (     a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     clk : in std_logic := '0';     sclr : IN STD_LOGIC;     ce : IN STD_LOGIC;     result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);     rdy : OUT STD_LOGIC   ); END Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692;  ARCHITECTURE Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692_a OF Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692 IS COMPONENT wrapped_Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692   PORT (     a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);     clk : IN STD_LOGIC;     sclr : IN STD_LOGIC;     ce : IN STD_LOGIC;     result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);     rdy : OUT STD_LOGIC   ); END COMPONENT;    FOR ALL : wrapped_Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692 USE ENTITY XilinxCoreLib.floating_point_v5_0(behavioral)     GENERIC MAP (       c_a_fraction_width => 24,       c_a_width => 32,       c_b_fraction_width => 24,       c_b_width => 32,       c_compare_operation => 8,       c_has_a_nd => 0,       c_has_a_negate => 0,       c_has_a_rfd => 0,       c_has_aclr => 0,       c_has_add => 0,       c_has_b_nd => 0,       c_has_b_negate => 0,       c_has_b_rfd => 0,       c_has_ce => 1,       c_has_compare => 0,       c_has_cts => 0,       c_has_divide => 0,       c_has_divide_by_zero => 0,       c_has_exception => 0,       c_has_fix_to_flt => 0,       c_has_flt_to_fix => 0,       c_has_flt_to_flt => 0,       c_has_inexact => 0,       c_has_invalid_op => 0,       c_has_multiply => 0,       c_has_operation_nd => 0,       c_has_operation_rfd => 0,       c_has_overflow => 0,       c_has_rdy => 1,       c_has_sclr => 1,       c_has_sqrt => 0,       c_has_status => 0,       c_has_subtract => 1,       c_has_underflow => 0,       c_latency => 1,       c_mult_usage => 0,       c_optimization => 1,       c_rate => 1,       c_result_fraction_width => 24,       c_result_width => 32,       c_speed => 2,       c_status_early => 0,       c_xdevicefamily => "spartan6"     ); BEGIN U0 : wrapped_Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692   PORT MAP (     a => a,     b => b,     clk => clk,     sclr => sclr,     ce => ce,     result => result,     rdy => rdy   );  END Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692_a; 
configuration conf_C3ADE5BE76064AA39E7EE6565DE88692 of Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692 is
  for Subtract_SCTL_L1_C3ADE5BE76064AA39E7EE6565DE88692_a end for; 
end conf_C3ADE5BE76064AA39E7EE6565DE88692; 