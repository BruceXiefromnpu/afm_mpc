  LIBRARY ieee; USE ieee.std_logic_1164.ALL; LIBRARY XilinxCoreLib; ENTITY Multiply_Accumulator_635C28D3DC43420AADC518895231A915 IS   PORT (     clk : in std_logic := '0';     ce : IN STD_LOGIC;     sclr : IN STD_LOGIC;     bypass : IN STD_LOGIC;     a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);     s : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)   ); END Multiply_Accumulator_635C28D3DC43420AADC518895231A915;  ARCHITECTURE Multiply_Accumulator_635C28D3DC43420AADC518895231A915_a OF Multiply_Accumulator_635C28D3DC43420AADC518895231A915 IS COMPONENT wrapped_Multiply_Accumulator_635C28D3DC43420AADC518895231A915   PORT (     clk : IN STD_LOGIC;     ce : IN STD_LOGIC;     sclr : IN STD_LOGIC;     bypass : IN STD_LOGIC;     a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);     b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);     s : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)   ); END COMPONENT;    FOR ALL : wrapped_Multiply_Accumulator_635C28D3DC43420AADC518895231A915 USE ENTITY XilinxCoreLib.xbip_multaccum_v2_0(behavioral)     GENERIC MAP (       c_a_type => 0,       c_a_width => 16,       c_accum_mode => 0,       c_accum_width => 32,       c_b_type => 0,       c_b_width => 16,       c_bypass_low => 0,       c_ce_overrides_sclr => 0,       c_has_bypass => 1,       c_latency => 1,       c_out_width => 32,       c_round_type => 0,       c_use_dsp48 => 1,       c_verbosity => 0,       c_xdevicefamily => "spartan6"     ); BEGIN U0 : wrapped_Multiply_Accumulator_635C28D3DC43420AADC518895231A915   PORT MAP (     clk => clk,     ce => ce,     sclr => sclr,     bypass => bypass,     a => a,     b => b,     s => s   );  END Multiply_Accumulator_635C28D3DC43420AADC518895231A915_a; 
configuration conf_635C28D3DC43420AADC518895231A915 of Multiply_Accumulator_635C28D3DC43420AADC518895231A915 is
  for Multiply_Accumulator_635C28D3DC43420AADC518895231A915_a end for; 
end conf_635C28D3DC43420AADC518895231A915; 